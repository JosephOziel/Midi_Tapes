BZh91AY&SY�/!h _�Py����߰����PrD��hR�� �`�2��� �`�2��H�(L�щ�6�	��� 4 E%jzj��� 4   �B�D�����Sjb2@���F��UF:�	�����D���Q�"""��|�@!�,��1]�Z86O�;����[�R�;&B��LQ����e�OLn%��R[M}eC6���L�$�
-�E�!�M{�[�]җ��f^aP�w�4��fϜL�eEo�P�~Q�/i�3fB���S�jD5� f��c�@��ge�͜r*�r���B��4��+���Pa��KeR�b̌�b�K��T]�h8զM���c��*S��W�a�""�Hw0��|"0�Yj@WI��R�,)`#$�F,�%Lߪ�a�ī��dB��X�1�k5Cndy�(P�%�h^U�՘��f�y�q�m���\�Cٝ_V�e;���K�J&aSF�,�O���,�A�JX*�8=�̩���M:\Z�r4{�[{�x�������xpM�)�ú��XY0��>d�;՗�H.��M�K��^!�u����5ׄ(Xt�(/�;�	Eß��*LV�t�ĚR�sq:���^���e����03Mp��Eo�H�jV�J���$J��I���L��A&¡�q�B���=�9i1�p���p�~`��� d!�H_�1`�=a�M{�-�E�^=t��w��G�w��O��)�9�e��	(�n`���X�r�a]
�	,���A�}}��#�#�?$!ł��Il� �ލ��`SX���Q���V$��AadT}5��E�/�b]��e/	B���s[�J�~S�Y��u=vұ]�v���NxP��*[�	���z����s	�<�iF$%����"���ሤ'g՟X�+���6�7!�7��(ؠ+ ��M�&��{'�iS���x�@�ߏぐ`�x��Z��N�ښ�çI�,���������F��'�P2׬�Б£�`@���fG�{D�/��2>�6�4ktx{ ��0C�Q� bt ^���H�
��- 